module hex_dump(
    input clk, rst, sig, fpga_rx,
    output fpga_tx, rdy3, rdy4,
);

    wire lock;
    assign rdy4 = value[3];
    assign rdy3 = sig;
    wire [7:0] value;
    dispatcher dispatcher(.clk(clk), .rst_in(rst), .sig(sig), .stb(stb), .value(value));

    reg tx_start;
    wire empty;
    wire full;
    wire [7:0] touart;
    fifo fifo(.clk(clk), .reset(rst), .wr(stb && !phase[0]), .rd(tx_start), .din(value), .empty(empty), .full(full), .dout(touart));
    reg [1:0] phase;
    reg [24:0] counter;

    always@(posedge clk)
    begin
        if (full) begin
            phase <= 1;
        end
        if ((!empty) && (!tx_busy) && (phase == 1)) begin
            tx_start <= 1;
        end else begin
            tx_start <= 0;
        end
        if (empty && (phase == 1)) begin
            phase <= 3;
        end
        if (phase == 3) begin
            counter <= counter - 1;
        end
        if ((phase == 3) && (counter == 0)) begin
            phase <= 0;
        end
    end

    wire tx_busy;
    localparam sym_rate = 1000000;
    localparam clk_freq = 48000000;
    localparam sym_cnt = clk_freq / sym_rate;
    localparam SCW = $clog2(sym_cnt);

    acia_tx #(
        .SCW(SCW),              // rate counter width
        .sym_cnt(sym_cnt)       // rate count value
    )
    my_tx(
        .clk(clk),				// system clock
        .rst(rst),			// system reset
        .tx_dat(touart),           // transmit data byte
        .tx_start(tx_start),    // trigger transmission
        .tx_serial(fpga_tx),         // tx serial output
        .tx_busy(tx_busy)       // tx is active (not ready)
    );

endmodule