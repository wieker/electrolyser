module top(
    output LED1, led2, led3
);

    assign LED1 = 1;
    assign led2 = 0;
    assign led3 = 1;

endmodule
