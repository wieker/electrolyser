module top(
    output LED1, LED2
);



    assign LED1 = 1;
    assign LED2 = 0;

endmodule
