module top(
    output LED1
);



    assign LED1 = 1;

endmodule
